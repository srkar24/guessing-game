library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity rand_gen_tb is

end rand_gen_tb;

architecture Behavioral of rand_gen_tb is

begin

end Behavioral;